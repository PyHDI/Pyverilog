//`default_nettype none

module TOP(CLK, RST);
  input CLK, RST;
  parameter AAA = 1;
  supply0 VSS;
  supply1 VDD;

endmodule

